module memory(
	input clk,

	// Control
	input d_read,
	input d_write,
	input d_push,
	input i_read,
	input i_push,

	// Buses
	input      [15:0] d_addr,
	input      [15:0] i_addr,
	inout      [15:0] d_bus
	);
	
	parameter mem_size = 512;

	(* ram_style = "block" *) reg [15:0] mem [mem_size-1:0];
	reg [15:0] m_store;
	assign d_bus = 
		i_push ? m_store :
		d_push ? m_store : 
		16'bz;

	integer i;
	initial begin
		for (i = 0; i < mem_size; i = i + 1) begin
			mem[i] = 16'b0;
		end

		//TODO: put default program here. Maybe it just displays hello world?
mem[0] = 16'b0000000000000000;
mem[1] = 16'b0000000000000000;
mem[2] = 16'b0000000000000000;
mem[3] = 16'b0000000000000000;
mem[4] = 16'b0000000000000000;
mem[5] = 16'b0000000000000000;
mem[6] = 16'b0000000000000000;
mem[7] = 16'b0000000000000000;
mem[8] = 16'b0000000000000000;
mem[9] = 16'b0000000000000000;
mem[10] = 16'b0000000000000000;
mem[11] = 16'b0000000000000000;
mem[12] = 16'b0000000000000000;
mem[13] = 16'b0000000000000000;
mem[14] = 16'b0000000000000000;
mem[15] = 16'b0000000000000000;
mem[16] = 16'b1011111100000001;
mem[17] = 16'b1100111100100011;
mem[18] = 16'b1011000000000000;
mem[19] = 16'b1100000000011000;
mem[20] = 16'b1111001111110000;
mem[21] = 16'b0000000000000000;
mem[22] = 16'b1111100101000000;
mem[23] = 16'b0000000000000000;
mem[24] = 16'b1011010100000000;
mem[25] = 16'b1100010100010110;
mem[26] = 16'b1011010000000000;
mem[27] = 16'b1100010000000000;
mem[28] = 16'b1111100101000000;
mem[29] = 16'b1011000000000000;
mem[30] = 16'b1100000000100101;
mem[31] = 16'b1011000100000000;
mem[32] = 16'b1100000100100101;
mem[33] = 16'b1111001000000001;
mem[34] = 16'b1111001101100101;
mem[35] = 16'b1011010000000000;
mem[36] = 16'b1100010000000001;
mem[37] = 16'b1111100101000000;
mem[38] = 16'b1011000000000000;
mem[39] = 16'b1100000000000111;
mem[40] = 16'b1011000100000000;
mem[41] = 16'b1100000100011101;
mem[42] = 16'b1011001100000000;
mem[43] = 16'b1100001100100100;
mem[44] = 16'b0001000000010010;
mem[45] = 16'b1111001000100011;
mem[46] = 16'b1111001101100101;
mem[47] = 16'b1011010000000000;
mem[48] = 16'b1100010000000010;
mem[49] = 16'b1111100101000000;
mem[50] = 16'b1011000000000000;
mem[51] = 16'b1100000000100100;
mem[52] = 16'b1011000100000000;
mem[53] = 16'b1100000100000111;
mem[54] = 16'b1011001100000000;
mem[55] = 16'b1100001100011101;
mem[56] = 16'b0010000000010010;
mem[57] = 16'b1111001000100011;
mem[58] = 16'b1111001101100101;
mem[59] = 16'b1011010000000000;
mem[60] = 16'b1100010000000011;
mem[61] = 16'b1111100101000000;
mem[62] = 16'b1011000000000000;
mem[63] = 16'b1100000000100100;
mem[64] = 16'b1011001100000000;
mem[65] = 16'b1100001100100101;
mem[66] = 16'b1111111100110000;
mem[67] = 16'b1111001000000011;
mem[68] = 16'b1111001101100101;
mem[69] = 16'b1011010000000000;
mem[70] = 16'b1100010000000100;
mem[71] = 16'b1111100101000000;
mem[72] = 16'b1011000000000000;
mem[73] = 16'b1100000000100100;
mem[74] = 16'b1011001100000000;
mem[75] = 16'b1100001100100011;
mem[76] = 16'b1111111101000000;
mem[77] = 16'b1111001000000011;
mem[78] = 16'b1111001101100101;
mem[79] = 16'b1011010000000000;
mem[80] = 16'b1100010000000110;
mem[81] = 16'b1111100101000000;
mem[82] = 16'b1011000000000000;
mem[83] = 16'b1100000000100100;
mem[84] = 16'b1011000100000000;
mem[85] = 16'b1100000100000111;
mem[86] = 16'b1011001100000000;
mem[87] = 16'b1100001111111100;
mem[88] = 16'b0011000000010010;
mem[89] = 16'b1111001000100011;
mem[90] = 16'b1111001101100101;
mem[91] = 16'b1011010000000000;
mem[92] = 16'b1100010000000111;
mem[93] = 16'b1111100101000000;
mem[94] = 16'b1011000000000000;
mem[95] = 16'b1100000000100100;
mem[96] = 16'b1011000100000000;
mem[97] = 16'b1100000100000111;
mem[98] = 16'b1011001100000000;
mem[99] = 16'b1100001100000101;
mem[100] = 16'b0100000000010010;
mem[101] = 16'b1111001000100011;
mem[102] = 16'b1111001101100101;
mem[103] = 16'b1011010000000000;
mem[104] = 16'b1100010000001000;
mem[105] = 16'b1111100101000000;
mem[106] = 16'b1011000000000000;
mem[107] = 16'b1100000000100100;
mem[108] = 16'b1011000100000000;
mem[109] = 16'b1100000100000111;
mem[110] = 16'b1011001100000000;
mem[111] = 16'b1100001100000001;
mem[112] = 16'b0101000000010010;
mem[113] = 16'b1111001000100011;
mem[114] = 16'b1111001101100101;
mem[115] = 16'b1011010000000000;
mem[116] = 16'b1100010000001001;
mem[117] = 16'b1111100101000000;
mem[118] = 16'b1011000000000000;
mem[119] = 16'b1100000000001000;
mem[120] = 16'b1011000100000000;
mem[121] = 16'b1100000100000010;
mem[122] = 16'b1011001100000000;
mem[123] = 16'b1100001100000010;
mem[124] = 16'b1001000000010010;
mem[125] = 16'b1111001000100011;
mem[126] = 16'b1111001101100101;
mem[127] = 16'b1011010000000000;
mem[128] = 16'b1100010000001010;
mem[129] = 16'b1111100101000000;
mem[130] = 16'b1011000000000000;
mem[131] = 16'b1100000000000010;
mem[132] = 16'b1011000100000000;
mem[133] = 16'b1100000100000011;
mem[134] = 16'b1011001100000000;
mem[135] = 16'b1100001100010000;
mem[136] = 16'b1010000000010010;
mem[137] = 16'b1111001000100011;
mem[138] = 16'b1011010000000000;
mem[139] = 16'b1100010000001011;
mem[140] = 16'b1111100101000000;
mem[141] = 16'b1011000000000000;
mem[142] = 16'b1100000000000101;
mem[143] = 16'b1011000100000000;
mem[144] = 16'b1100000100000110;
mem[145] = 16'b1011001100000000;
mem[146] = 16'b1100001100000100;
mem[147] = 16'b0110000000010010;
mem[148] = 16'b1111001000100011;
mem[149] = 16'b1111001101100101;
mem[150] = 16'b1011010000000000;
mem[151] = 16'b1100010000001100;
mem[152] = 16'b1111100101000000;
mem[153] = 16'b1011000000000000;
mem[154] = 16'b1100000000000101;
mem[155] = 16'b1011000100000000;
mem[156] = 16'b1100000100000110;
mem[157] = 16'b1011001100000000;
mem[158] = 16'b1100001100000111;
mem[159] = 16'b0111000000010010;
mem[160] = 16'b1111001000100011;
mem[161] = 16'b1111001101100101;
mem[162] = 16'b1011010000000000;
mem[163] = 16'b1100010000001101;
mem[164] = 16'b1111100101000000;
mem[165] = 16'b1011000000000000;
mem[166] = 16'b1100000000000101;
mem[167] = 16'b1011000100000000;
mem[168] = 16'b1100000100000110;
mem[169] = 16'b1011001100000000;
mem[170] = 16'b1100001100000011;
mem[171] = 16'b1000000000010010;
mem[172] = 16'b1111001000100011;
mem[173] = 16'b1111001101100101;
mem[174] = 16'b1011010000000000;
mem[175] = 16'b1100010000001110;
mem[176] = 16'b1111100101000000;
mem[177] = 16'b1011000000000100;
mem[178] = 16'b1100000011110011;
mem[179] = 16'b1011001111111011;
mem[180] = 16'b1100001100001100;
mem[181] = 16'b1111011000000010;
mem[182] = 16'b1111001000100011;
mem[183] = 16'b1111001101100101;
mem[184] = 16'b1011010000000000;
mem[185] = 16'b1100010000001111;
mem[186] = 16'b1111100101000000;
mem[187] = 16'b1011000000000100;
mem[188] = 16'b1100000011110011;
mem[189] = 16'b1011001100000100;
mem[190] = 16'b1100001111110011;
mem[191] = 16'b1111000100000010;
mem[192] = 16'b1111001000100011;
mem[193] = 16'b1111001101100101;
mem[194] = 16'b1011010000000000;
mem[195] = 16'b1100010000010000;
mem[196] = 16'b1111100101000000;
mem[197] = 16'b1011000000000000;
mem[198] = 16'b1100000000001010;
mem[199] = 16'b1111000111110001;
mem[200] = 16'b1111101000001111;
mem[201] = 16'b1111111100110001;
mem[202] = 16'b1111001000011111;
mem[203] = 16'b1111001101100101;
mem[204] = 16'b1111111101000001;
mem[205] = 16'b1111010000010010;
mem[206] = 16'b1111001000000010;
mem[207] = 16'b1111001101100101;
mem[208] = 16'b1011010000000000;
mem[209] = 16'b1100010000010001;
mem[210] = 16'b1111100101000000;
mem[211] = 16'b1011000000000000;
mem[212] = 16'b1100000000001100;
mem[213] = 16'b1111000111110001;
mem[214] = 16'b1111101000001111;
mem[215] = 16'b1111101111110010;
mem[216] = 16'b1111001000011111;
mem[217] = 16'b1111001101100101;
mem[218] = 16'b1111001000000010;
mem[219] = 16'b1111001101100101;
mem[220] = 16'b1011010000000000;
mem[221] = 16'b1100010000010010;
mem[222] = 16'b1111100101000000;
mem[223] = 16'b1011000000000001;
mem[224] = 16'b1100000000100001;
mem[225] = 16'b1011001100000000;
mem[226] = 16'b1100001101111111;
mem[227] = 16'b1111010000000010;
mem[228] = 16'b1111001000100011;
mem[229] = 16'b1111001101100101;
mem[230] = 16'b1011010000000000;
mem[231] = 16'b1100010000010011;
mem[232] = 16'b1111100101000000;
mem[233] = 16'b1011000000000001;
mem[234] = 16'b1100000000100001;
mem[235] = 16'b1011001100000000;
mem[236] = 16'b1100001101001100;
mem[237] = 16'b1111010100110000;
mem[238] = 16'b1111010000000010;
mem[239] = 16'b1111001000100011;
mem[240] = 16'b1111001101100101;
mem[241] = 16'b1011010000000000;
mem[242] = 16'b1100010000010100;
mem[243] = 16'b1111100101000000;
mem[244] = 16'b1011000000000000;
mem[245] = 16'b1100000001001001;
mem[246] = 16'b1011001100000000;
mem[247] = 16'b1100001101001001;
mem[248] = 16'b1111100100000000;
mem[249] = 16'b1111100000000010;
mem[250] = 16'b1011000000000000;
mem[251] = 16'b1100000000000000;
mem[252] = 16'b1111100100000000;
mem[253] = 16'b1111001000100011;
mem[254] = 16'b1111001101100101;
mem[255] = 16'b1011010000000000;
mem[256] = 16'b1100010000010101;
mem[257] = 16'b1111100101000000;
mem[258] = 16'b1011000000000000;
mem[259] = 16'b1100000000000101;
mem[260] = 16'b1111001000000100;
mem[261] = 16'b1111111100100000;
mem[262] = 16'b1111001101100101;
mem[263] = 16'b1011010000000000;
mem[264] = 16'b1100010000010110;
mem[265] = 16'b1111100101000000;
mem[266] = 16'b1011000000000000;
mem[267] = 16'b1100000000000100;
mem[268] = 16'b1011001100000000;
mem[269] = 16'b1100001100000100;
mem[270] = 16'b1111111100100000;
mem[271] = 16'b1111111100010010;
mem[272] = 16'b1111001000100011;
mem[273] = 16'b1111001101100101;
mem[274] = 16'b1011010000000000;
mem[275] = 16'b1100010000010111;
mem[276] = 16'b1111100101000000;
mem[277] = 16'b1011000000000001;
mem[278] = 16'b1100000000011011;
mem[279] = 16'b1011001100000001;
mem[280] = 16'b1100001100011010;
mem[281] = 16'b1111110000000010;
mem[282] = 16'b1111001111110101;
mem[283] = 16'b1111001000100011;
mem[284] = 16'b1111001101100101;
mem[285] = 16'b1011000000000000;
mem[286] = 16'b1100000011111111;
mem[287] = 16'b1111100100000000;
mem[288] = 16'b0000000000000000;
mem[289] = 16'b0000000001111111;
mem[290] = 16'b0000000000000000;


	end
	
	assign read = d_read || i_read;
	wire [15:0] addr;
	assign addr = 
		d_read ? d_addr :
		i_read ? i_addr :
		d_addr;

	always @ (posedge clk) begin
		if (read) begin
			m_store <= mem[addr];
		end else if (d_write) begin
			mem[addr] <= d_bus;
		end
	end

endmodule
