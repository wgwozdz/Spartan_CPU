module memory(
	input clk,

	// Control
	input d_read,
	input d_write,
	input d_push,
	input i_read,
	input i_push,

	// Buses
	input      [15:0] d_addr,
	input      [15:0] i_addr,
	inout      [15:0] d_bus
	);

	(* ram_style = "block" *) reg [15:0] mem [255:0];
	reg [15:0] m_store;
	assign d_bus = 
		i_push ? m_store :
		d_push ? m_store : 
		16'bz;

	integer i;
	initial begin
		for (i = 0; i < 256; i = i + 1) begin
			mem[i] = 16'b0;
		end

		//TODO: put default program here. Maybe it just displays hello world?

mem[0] = 16'b0000000000000000;
mem[1] = 16'b0000000000000000;
mem[2] = 16'b0000000000000000;
mem[3] = 16'b0000000000000000;
mem[4] = 16'b0000000000000000;
mem[5] = 16'b0000000000000000;
mem[6] = 16'b0000000000000000;
mem[7] = 16'b0000000000000000;
mem[8] = 16'b0000000000000000;
mem[9] = 16'b0000000000000000;
mem[10] = 16'b0000000000000000;
mem[11] = 16'b0000000000000000;
mem[12] = 16'b0000000000000000;
mem[13] = 16'b0000000000000000;
mem[14] = 16'b0000000000000000;
mem[15] = 16'b0000000000000000;
mem[16] = 16'b1011111100000000;
mem[17] = 16'b1100111110110000;
mem[18] = 16'b1011000000000000;
mem[19] = 16'b1100000000011000;
mem[20] = 16'b1111001101110000;
mem[21] = 16'b0000000000000000;
mem[22] = 16'b1111100101000000;
mem[23] = 16'b0000000000000000;
mem[24] = 16'b1011010100000000;
mem[25] = 16'b1100010100010110;
mem[26] = 16'b1011010000000000;
mem[27] = 16'b1100010000000000;
mem[28] = 16'b1011000000000000;
mem[29] = 16'b1100000000100101;
mem[30] = 16'b1011000100000000;
mem[31] = 16'b1100000100100101;
mem[32] = 16'b1111001000000001;
mem[33] = 16'b1111001101100101;
mem[34] = 16'b1011010000000000;
mem[35] = 16'b1100010000000001;
mem[36] = 16'b1011000000000000;
mem[37] = 16'b1100000000000111;
mem[38] = 16'b1011000100000000;
mem[39] = 16'b1100000100011101;
mem[40] = 16'b1011001100000000;
mem[41] = 16'b1100001100100100;
mem[42] = 16'b0001000000010010;
mem[43] = 16'b1111001000100011;
mem[44] = 16'b1111001101100101;
mem[45] = 16'b1011010000000000;
mem[46] = 16'b1100010000000010;
mem[47] = 16'b1011000000000000;
mem[48] = 16'b1100000000100100;
mem[49] = 16'b1011000100000000;
mem[50] = 16'b1100000100000111;
mem[51] = 16'b1011001100000000;
mem[52] = 16'b1100001100011101;
mem[53] = 16'b0010000000010010;
mem[54] = 16'b1111001000100011;
mem[55] = 16'b1111001101100101;
mem[56] = 16'b1011010000000000;
mem[57] = 16'b1100010000000011;
mem[58] = 16'b1011000000000000;
mem[59] = 16'b1100000000100100;
mem[60] = 16'b1011001100000000;
mem[61] = 16'b1100001100100101;
mem[62] = 16'b1111111100110000;
mem[63] = 16'b1111001000000011;
mem[64] = 16'b1111001101100101;
mem[65] = 16'b1011010000000000;
mem[66] = 16'b1100010000000100;
mem[67] = 16'b1011000000000000;
mem[68] = 16'b1100000000100100;
mem[69] = 16'b1011001100000000;
mem[70] = 16'b1100001100100011;
mem[71] = 16'b1111111101000000;
mem[72] = 16'b1111001000000011;
mem[73] = 16'b1111001101100101;
mem[74] = 16'b1011010000000000;
mem[75] = 16'b1100010000000110;
mem[76] = 16'b1011000000000000;
mem[77] = 16'b1100000000100100;
mem[78] = 16'b1011000100000000;
mem[79] = 16'b1100000100000111;
mem[80] = 16'b1011001100000000;
mem[81] = 16'b1100001111111100;
mem[82] = 16'b0011000000010010;
mem[83] = 16'b1111001000100011;
mem[84] = 16'b1111001101100101;
mem[85] = 16'b1011010000000000;
mem[86] = 16'b1100010000000111;
mem[87] = 16'b1011000000000000;
mem[88] = 16'b1100000000100100;
mem[89] = 16'b1011000100000000;
mem[90] = 16'b1100000100000111;
mem[91] = 16'b1011001100000000;
mem[92] = 16'b1100001100000101;
mem[93] = 16'b0100000000010010;
mem[94] = 16'b1111001000100011;
mem[95] = 16'b1111001101100101;
mem[96] = 16'b1011010000000000;
mem[97] = 16'b1100010000001000;
mem[98] = 16'b1011000000000000;
mem[99] = 16'b1100000000100100;
mem[100] = 16'b1011000100000000;
mem[101] = 16'b1100000100000111;
mem[102] = 16'b1011001100000000;
mem[103] = 16'b1100001100000001;
mem[104] = 16'b0101000000010010;
mem[105] = 16'b1111001000100011;
mem[106] = 16'b1111001101100101;
mem[107] = 16'b1011010000000000;
mem[108] = 16'b1100010000001001;
mem[109] = 16'b1011000000000000;
mem[110] = 16'b1100000000001000;
mem[111] = 16'b1011000100000000;
mem[112] = 16'b1100000100000010;
mem[113] = 16'b1011001100000000;
mem[114] = 16'b1100001100000010;
mem[115] = 16'b1001000000010010;
mem[116] = 16'b1111001000100011;
mem[117] = 16'b1111001101100101;
mem[118] = 16'b1011010000000000;
mem[119] = 16'b1100010000001010;
mem[120] = 16'b1011000000000000;
mem[121] = 16'b1100000000000010;
mem[122] = 16'b1011000100000000;
mem[123] = 16'b1100000100000011;
mem[124] = 16'b1011001100000000;
mem[125] = 16'b1100001100010000;
mem[126] = 16'b1010000000010010;
mem[127] = 16'b1111001000100011;
mem[128] = 16'b1111001101100101;
mem[129] = 16'b1011010000000000;
mem[130] = 16'b1100010000001011;
mem[131] = 16'b1011000000000000;
mem[132] = 16'b1100000000000101;
mem[133] = 16'b1011000100000000;
mem[134] = 16'b1100000100000110;
mem[135] = 16'b1011001100000000;
mem[136] = 16'b1100001100000100;
mem[137] = 16'b0110000000010010;
mem[138] = 16'b1111001000100011;
mem[139] = 16'b1111001101100101;
mem[140] = 16'b1011010000000000;
mem[141] = 16'b1100010000001100;
mem[142] = 16'b1011000000000000;
mem[143] = 16'b1100000000000101;
mem[144] = 16'b1011000100000000;
mem[145] = 16'b1100000100000110;
mem[146] = 16'b1011001100000000;
mem[147] = 16'b1100001100000111;
mem[148] = 16'b0111000000010010;
mem[149] = 16'b1111001000100011;
mem[150] = 16'b1111001101100101;
mem[151] = 16'b1011010000000000;
mem[152] = 16'b1100010000001101;
mem[153] = 16'b1011000000000000;
mem[154] = 16'b1100000000000101;
mem[155] = 16'b1011000100000000;
mem[156] = 16'b1100000100000110;
mem[157] = 16'b1011001100000000;
mem[158] = 16'b1100001100000011;
mem[159] = 16'b1000000000010010;
mem[160] = 16'b1111001000100011;
mem[161] = 16'b1111001101100101;
mem[162] = 16'b1011010000000000;
mem[163] = 16'b1100010000001110;
mem[164] = 16'b1011000000000100;
mem[165] = 16'b1100000011110011;
mem[166] = 16'b1011001111111011;
mem[167] = 16'b1100001100001100;
mem[168] = 16'b1111011000000010;
mem[169] = 16'b1111001000100011;
mem[170] = 16'b1111001101100101;
mem[171] = 16'b1011000000000000;
mem[172] = 16'b1100000011111111;
mem[173] = 16'b1111100100000000;
mem[174] = 16'b0000000000000000;
mem[175] = 16'b0000000000000000;



	end
	
	assign read = d_read || i_read;
	wire [15:0] addr;
	assign addr = 
		d_read ? d_addr :
		i_read ? i_addr :
		d_addr;

	always @ (posedge clk) begin
		if (read) begin
			m_store <= mem[addr];
		end else if (d_write) begin
			mem[addr] <= d_bus;
		end
	end

endmodule
